module Datapath();
endmodule